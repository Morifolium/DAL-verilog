module new_fp16_add_timing (
    
);
    
endmodule