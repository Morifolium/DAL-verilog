// Copyright 2019 ETH Zurich and University of Bologna.
//
// Copyright and related rights are licensed under the Solderpad Hardware
// License, Version 0.51 (the "License"); you may not use this file except in
// compliance with the License. You may obtain a copy of the License at
// http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
// or agreed to in writing, software, hardware and materials distributed under
// this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
// CONDITIONS OF ANY KIND, either express or implied. See the License for the
// specific language governing permissions and limitations under the License.
//
// SPDX-License-Identifier: SHL-0.51

// Author: Stefan Mach <smach@iis.ee.ethz.ch>


module fpnew_classifier #(
    parameter  fpnew_pkg::fp_format_e FpFormat    = fpnew_pkg::fp_format_e'(2),
    parameter  int unsigned           NumOperands = 1,
    // Do not change
    localparam int unsigned           WIDTH       = fpnew_pkg::fp_width(FpFormat)
) (
    input  logic                [NumOperands-1:0][WIDTH-1:0] operands_i,
    input  logic                [NumOperands-1:0]            is_boxed_i,
    output fpnew_pkg::fp_info_t [NumOperands-1:0]            info_o
);

  localparam int unsigned EXP_BITS = fpnew_pkg::exp_bits(FpFormat);
  localparam int unsigned MAN_BITS = fpnew_pkg::man_bits(FpFormat);

  // Type definition
  typedef struct packed {
    logic                sign;
    logic [EXP_BITS-1:0] exponent;
    logic [MAN_BITS-1:0] mantissa;
  } fp_t;

  // Iterate through all operands
  for (genvar op = 0; op < int'(NumOperands); op++) begin : gen_num_values

    fp_t  value;
    logic is_boxed;
    logic is_normal;
    logic is_inf;
    logic is_nan;
    logic is_signalling;
    logic is_quiet;
    logic is_zero;
    logic is_subnormal;

    // ---------------
    // Classify Input
    // ---------------
    //only consider  normal/subnormal/zero
    always_comb begin : classify_input
      value                    = operands_i[op];
      //is_boxed      = is_boxed_i[op];
      is_boxed                 = 1'b1;
      is_normal                = is_boxed && (value.exponent != '0) && (value.exponent != '1);
      is_zero                  = is_boxed && (value.exponent == '0) && (value.mantissa == '0);
      is_subnormal             = is_boxed && (value.exponent == '0) && !is_zero;

      //is_inf        = is_boxed && ((value.exponent == '1) && (value.mantissa == '0));
      is_inf                   = 1'b0;
      //is_nan        = !is_boxed || ((value.exponent == '1) && (value.mantissa != '0));
      is_nan                   = 1'b0;
      //is_signalling = is_boxed && is_nan && (value.mantissa[MAN_BITS-1] == 1'b0);
      is_signalling            = 1'b0;
      //is_quiet                 = is_nan && !is_signalling;
      is_quiet                 = 1'b0;
      // Assign output for current input
      info_o[op].is_normal     = is_normal;
      info_o[op].is_subnormal  = is_subnormal;
      info_o[op].is_zero       = is_zero;
      info_o[op].is_inf        = is_inf;
      info_o[op].is_nan        = is_nan;
      info_o[op].is_signalling = is_signalling;
      info_o[op].is_quiet      = is_quiet;
      info_o[op].is_boxed      = is_boxed;
    end




  end
endmodule
